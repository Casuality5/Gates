module NOT(
    input wire a,
    output wire y
);
    assign y=~a;
endmodule